`define REGREAD_SECURE
`define REGWRITE_SECURE
`define MEM_SECURE
`define RV_A 3
`define RV_B 2
//`define MD_SECURE
`define SHIFT_SECURE
`define ADDER_SECURE
//`define CSR_SECURE